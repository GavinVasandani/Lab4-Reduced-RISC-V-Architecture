//Creating mux that's after regFile